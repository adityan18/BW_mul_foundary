`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 30.04.2022 15:52:18
// Design Name:
// Module Name: RAM
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module ram2
    #(
         //parameter ADDR_WIDTH = 10,
         parameter ADDR_WIDTH = 12,
         parameter MAX_FEATURES = 15,
         parameter LENGTH = 16,      //Num_data points
         parameter DATA_WIDTH = LENGTH * (MAX_FEATURES+1), //width = num_features + 1 for y values
         parameter DEPTH = 100     //Num_data points
         // parameter DEPTH = 4      //Num_data points
         //parameter LEN_BITS = 4     // Num_bits required to get 'LENGTH' features
     )
     (
         input oe, we, RST,
         input [ADDR_WIDTH-1:0] addr,
         inout [DATA_WIDTH-1:0] data
     );
    //512kb

    integer i;
    reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];
    reg [DATA_WIDTH-1:0] buffer;
    //4 bits for features, 10 bits for data points

    //For Writing, enable cs, we, and make sure data is available at data bus on posedge.
    always@(addr or RST or we)
    begin
        if(RST)
        begin
            for(i=0;i<DEPTH;i=i+1)
            begin
                mem[i]<=0;
            end
        end
        else if(we)
        begin
            $display("%h", data);
            mem[addr] <= data;
        end
    end

    //For Reading, enable cs, oe, disable we, and data will be available on data bus at posedge
    always@(addr)
    begin
        if(~we)
        begin
            buffer <= mem[addr];
        end
    end

    assign data = (~we && oe) ? buffer : 'hz;

endmodule
