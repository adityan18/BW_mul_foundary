VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END a[0]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 0.000 421.730 4.000 ;
    END
  END a[7]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 0.000 477.850 4.000 ;
    END
  END b[0]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 0.000 533.970 4.000 ;
    END
  END b[1]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END b[2]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 0.000 702.330 4.000 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 0.000 758.450 4.000 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 0.000 814.570 4.000 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 0.000 870.690 4.000 ;
    END
  END b[7]
  PIN p[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 596.000 56.950 600.000 ;
    END
  END p[0]
  PIN p[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 596.000 169.190 600.000 ;
    END
  END p[1]
  PIN p[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 596.000 281.430 600.000 ;
    END
  END p[2]
  PIN p[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 596.000 393.670 600.000 ;
    END
  END p[3]
  PIN p[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 596.000 505.910 600.000 ;
    END
  END p[4]
  PIN p[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 596.000 618.150 600.000 ;
    END
  END p[5]
  PIN p[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 596.000 730.390 600.000 ;
    END
  END p[6]
  PIN p[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.350 596.000 842.630 600.000 ;
    END
  END p[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 583.385 894.430 586.215 ;
        RECT 5.330 577.945 894.430 580.775 ;
        RECT 5.330 572.505 894.430 575.335 ;
        RECT 5.330 567.065 894.430 569.895 ;
        RECT 5.330 561.625 894.430 564.455 ;
        RECT 5.330 556.185 894.430 559.015 ;
        RECT 5.330 550.745 894.430 553.575 ;
        RECT 5.330 545.305 894.430 548.135 ;
        RECT 5.330 539.865 894.430 542.695 ;
        RECT 5.330 534.425 894.430 537.255 ;
        RECT 5.330 528.985 894.430 531.815 ;
        RECT 5.330 523.545 894.430 526.375 ;
        RECT 5.330 518.105 894.430 520.935 ;
        RECT 5.330 512.665 894.430 515.495 ;
        RECT 5.330 507.225 894.430 510.055 ;
        RECT 5.330 501.785 894.430 504.615 ;
        RECT 5.330 496.345 894.430 499.175 ;
        RECT 5.330 490.905 894.430 493.735 ;
        RECT 5.330 485.465 894.430 488.295 ;
        RECT 5.330 480.025 894.430 482.855 ;
        RECT 5.330 474.585 894.430 477.415 ;
        RECT 5.330 469.145 894.430 471.975 ;
        RECT 5.330 463.705 894.430 466.535 ;
        RECT 5.330 458.265 894.430 461.095 ;
        RECT 5.330 452.825 894.430 455.655 ;
        RECT 5.330 447.385 894.430 450.215 ;
        RECT 5.330 441.945 894.430 444.775 ;
        RECT 5.330 436.505 894.430 439.335 ;
        RECT 5.330 431.065 894.430 433.895 ;
        RECT 5.330 425.625 894.430 428.455 ;
        RECT 5.330 420.185 894.430 423.015 ;
        RECT 5.330 414.745 894.430 417.575 ;
        RECT 5.330 409.305 894.430 412.135 ;
        RECT 5.330 403.865 894.430 406.695 ;
        RECT 5.330 398.425 894.430 401.255 ;
        RECT 5.330 392.985 894.430 395.815 ;
        RECT 5.330 387.545 894.430 390.375 ;
        RECT 5.330 382.105 894.430 384.935 ;
        RECT 5.330 376.665 894.430 379.495 ;
        RECT 5.330 371.225 894.430 374.055 ;
        RECT 5.330 365.785 894.430 368.615 ;
        RECT 5.330 360.345 894.430 363.175 ;
        RECT 5.330 354.905 894.430 357.735 ;
        RECT 5.330 349.465 894.430 352.295 ;
        RECT 5.330 344.025 894.430 346.855 ;
        RECT 5.330 338.585 894.430 341.415 ;
        RECT 5.330 333.145 894.430 335.975 ;
        RECT 5.330 327.705 894.430 330.535 ;
        RECT 5.330 322.265 894.430 325.095 ;
        RECT 5.330 316.825 894.430 319.655 ;
        RECT 5.330 311.385 894.430 314.215 ;
        RECT 5.330 305.945 894.430 308.775 ;
        RECT 5.330 300.505 894.430 303.335 ;
        RECT 5.330 295.065 894.430 297.895 ;
        RECT 5.330 289.625 894.430 292.455 ;
        RECT 5.330 284.185 894.430 287.015 ;
        RECT 5.330 278.745 894.430 281.575 ;
        RECT 5.330 273.305 894.430 276.135 ;
        RECT 5.330 267.865 894.430 270.695 ;
        RECT 5.330 262.425 894.430 265.255 ;
        RECT 5.330 256.985 894.430 259.815 ;
        RECT 5.330 251.545 894.430 254.375 ;
        RECT 5.330 246.105 894.430 248.935 ;
        RECT 5.330 240.665 894.430 243.495 ;
        RECT 5.330 235.225 894.430 238.055 ;
        RECT 5.330 229.785 894.430 232.615 ;
        RECT 5.330 224.345 894.430 227.175 ;
        RECT 5.330 218.905 894.430 221.735 ;
        RECT 5.330 213.465 894.430 216.295 ;
        RECT 5.330 208.025 894.430 210.855 ;
        RECT 5.330 202.585 894.430 205.415 ;
        RECT 5.330 197.145 894.430 199.975 ;
        RECT 5.330 191.705 894.430 194.535 ;
        RECT 5.330 186.265 894.430 189.095 ;
        RECT 5.330 180.825 894.430 183.655 ;
        RECT 5.330 175.385 894.430 178.215 ;
        RECT 5.330 169.945 894.430 172.775 ;
        RECT 5.330 164.505 894.430 167.335 ;
        RECT 5.330 159.065 894.430 161.895 ;
        RECT 5.330 153.625 894.430 156.455 ;
        RECT 5.330 148.185 894.430 151.015 ;
        RECT 5.330 142.745 894.430 145.575 ;
        RECT 5.330 137.305 894.430 140.135 ;
        RECT 5.330 131.865 894.430 134.695 ;
        RECT 5.330 126.425 894.430 129.255 ;
        RECT 5.330 120.985 894.430 123.815 ;
        RECT 5.330 115.545 894.430 118.375 ;
        RECT 5.330 110.105 894.430 112.935 ;
        RECT 5.330 104.665 894.430 107.495 ;
        RECT 5.330 99.225 894.430 102.055 ;
        RECT 5.330 93.785 894.430 96.615 ;
        RECT 5.330 88.345 894.430 91.175 ;
        RECT 5.330 82.905 894.430 85.735 ;
        RECT 5.330 77.465 894.430 80.295 ;
        RECT 5.330 72.025 894.430 74.855 ;
        RECT 5.330 66.585 894.430 69.415 ;
        RECT 5.330 61.145 894.430 63.975 ;
        RECT 5.330 55.705 894.430 58.535 ;
        RECT 5.330 50.265 894.430 53.095 ;
        RECT 5.330 44.825 894.430 47.655 ;
        RECT 5.330 39.385 894.430 42.215 ;
        RECT 5.330 33.945 894.430 36.775 ;
        RECT 5.330 28.505 894.430 31.335 ;
        RECT 5.330 23.065 894.430 25.895 ;
        RECT 5.330 17.625 894.430 20.455 ;
        RECT 5.330 12.185 894.430 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 9.220 894.240 587.760 ;
      LAYER met2 ;
        RECT 21.070 595.720 56.390 596.770 ;
        RECT 57.230 595.720 168.630 596.770 ;
        RECT 169.470 595.720 280.870 596.770 ;
        RECT 281.710 595.720 393.110 596.770 ;
        RECT 393.950 595.720 505.350 596.770 ;
        RECT 506.190 595.720 617.590 596.770 ;
        RECT 618.430 595.720 729.830 596.770 ;
        RECT 730.670 595.720 842.070 596.770 ;
        RECT 842.910 595.720 872.060 596.770 ;
        RECT 21.070 4.280 872.060 595.720 ;
        RECT 21.070 4.000 28.330 4.280 ;
        RECT 29.170 4.000 84.450 4.280 ;
        RECT 85.290 4.000 140.570 4.280 ;
        RECT 141.410 4.000 196.690 4.280 ;
        RECT 197.530 4.000 252.810 4.280 ;
        RECT 253.650 4.000 308.930 4.280 ;
        RECT 309.770 4.000 365.050 4.280 ;
        RECT 365.890 4.000 421.170 4.280 ;
        RECT 422.010 4.000 477.290 4.280 ;
        RECT 478.130 4.000 533.410 4.280 ;
        RECT 534.250 4.000 589.530 4.280 ;
        RECT 590.370 4.000 645.650 4.280 ;
        RECT 646.490 4.000 701.770 4.280 ;
        RECT 702.610 4.000 757.890 4.280 ;
        RECT 758.730 4.000 814.010 4.280 ;
        RECT 814.850 4.000 870.130 4.280 ;
        RECT 870.970 4.000 872.060 4.280 ;
      LAYER met3 ;
        RECT 21.050 10.715 867.430 587.685 ;
  END
END user_proj_example
END LIBRARY

